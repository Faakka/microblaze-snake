`timescale 1ns / 1ps

module hdmi_ctrl_tb;



endmodule
